`timescale 1ns / 1ps

module FSM(
input clk,
input rst,
input forward,
output state
    );
    



endmodule
